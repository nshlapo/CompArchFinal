module fp_adder
(
  input[31:0] A, B,
  output[31:0] Out
);

endmodule
