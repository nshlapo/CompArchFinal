module sqrt
(
  input[31:0] A,
  input sqrt_clk
  input fp_clk,
  input int_clk,
  output[31:0] Out
);

endmodule
