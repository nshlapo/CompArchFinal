module fp_divider
(
  input[31:0] A, B,
  input fp_clk,
  input int_clk,
  output[31:0] Out
);

endmodule
